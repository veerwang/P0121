	module main;

initial
begin
	$display("Hello world");
	$finish;
end

endmodule
